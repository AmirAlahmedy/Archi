
Library IEEE;
USE IEEE.std_logic_1164.all;
Entity DecALUREG is

  Port(clk,rst: in std_logic; 
Rdst :in std_logic_vector(15 downto 0);
 Rsrc: in std_logic_vector(15 downto 0);
Rdstout :out std_logic_vector(15 downto 0);
 Rsrcout: out std_logic_vector(15 downto 0);
Atype:in std_logic;
Aluop:in std_logic;
RegWrite:in std_logic;
Atypeout:out std_logic;
Aluopout:out std_logic;
RegWriteout:out std_logic;
RdstAddress : out std_logic_vector (2 downto 0);
RdstAddressIn : in std_logic_vector (2 downto 0);
shamtin:in std_logic_vector(4 downto 0);
shamtout:out std_logic_vector(4 downto 0);
Funcin:in std_logic_vector(2 downto 0);
funcout:out std_logic_vector(2 downto 0)

);
  end DecALUREG;
  
  architecture a_FetDecReg of DecALUREG is 
  begin
    process(clk)
      begin
        if(rst='1') then
funcout<="000";
shamtout<="00000";
Atypeout<='0';
Aluopout<='0';
RegWriteout<='0';
RdstAddress<="000";
      Rdstout<= (others=>'0');
 Rsrcout<= (others=>'0');
      elsif rising_edge(clk) then
shamtout<=shamtin;
Atypeout<=Atype;
Aluopout<=Aluop;
RegWriteout<=rEGwRITE;
    Rdstout<= Rdst;
RdstAddress<=RdstAddressIn;
 Rsrcout<= Rsrc;
funcout<=funcin;
      end if;
    end process;
   end ARCHITECTURE;